library verilog;
use verilog.vl_types.all;
entity cpu_test_sim_vlg_vec_tst is
end cpu_test_sim_vlg_vec_tst;
