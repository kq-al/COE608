library verilog;
use verilog.vl_types.all;
entity adder1_vlg_vec_tst is
end adder1_vlg_vec_tst;
