library verilog;
use verilog.vl_types.all;
entity alu32_vlg_vec_tst is
end alu32_vlg_vec_tst;
